`include "parameters.svh"

module wave_table_sine
    (
	    input reg [DATA_WIDTH-1:0] phase,
        output reg signed [DATA_WIDTH-1:0] signal
    );

    reg [DATA_WIDTH-1:0] sine_table [0:SINE_RESOLUTION-1] = {2047,2057,2068,2079,2089,2100,2111,2122,2132,2143,2154,2164,2175,2186,2196,2207,2218,2228,2239,2250,2260,2271,2282,2292,2303,2314,2324,2335,2346,2356,2367,2377,2388,2398,2409,2420,2430,2441,2451,2462,2472,2483,2493,2503,2514,2524,2535,2545,2556,2566,2576,2587,2597,2607,2618,2628,2638,2648,2659,2669,2679,2689,2699,2710,2720,2730,2740,2750,2760,2770,2780,2790,2800,2810,2820,2830,2840,2850,2859,2869,2879,2889,2899,2908,2918,2928,2937,2947,2957,2966,2976,2985,2995,3004,3014,3023,3033,3042,3051,3061,3070,3079,3089,3098,3107,3116,3125,3134,3143,3152,3161,3170,3179,3188,3197,3206,3215,3224,3232,3241,3250,3258,3267,3276,3284,3293,3301,3310,3318,3326,3335,3343,3351,3360,3368,3376,3384,3392,3400,3408,3416,3424,3432,3440,3448,3456,3463,3471,3479,3486,3494,3502,3509,3517,3524,3531,3539,3546,3553,3561,3568,3575,3582,3589,3596,3603,3610,3617,3624,3631,3637,3644,3651,3657,3664,3670,3677,3683,3690,3696,3703,3709,3715,3721,3727,3733,3740,3746,3751,3757,3763,3769,3775,3781,3786,3792,3797,3803,3808,3814,3819,3825,3830,3835,3840,3845,3851,3856,3861,3865,3870,3875,3880,3885,3889,3894,3899,3903,3908,3912,3917,3921,3925,3929,3934,3938,3942,3946,3950,3954,3958,3961,3965,3969,3972,3976,3980,3983,3987,3990,3993,3997,4000,4003,4006,4009,4012,4015,4018,4021,4024,4026,4029,4032,4034,4037,4039,4042,4044,4047,4049,4051,4053,4055,4057,4059,4061,4063,4065,4067,4068,4070,4072,4073,4075,4076,4077,4079,4080,4081,4082,4083,4084,4085,4086,4087,4088,4089,4089,4090,4091,4091,4092,4092,4092,4093,4093,4093,4093,4093,4094,4093,4093,4093,4093,4093,4092,4092,4092,4091,4091,4090,4089,4089,4088,4087,4086,4085,4084,4083,4082,4081,4080,4079,4077,4076,4075,4073,4072,4070,4068,4067,4065,4063,4061,4059,4057,4055,4053,4051,4049,4047,4044,4042,4039,4037,4034,4032,4029,4026,4024,4021,4018,4015,4012,4009,4006,4003,4000,3997,3993,3990,3987,3983,3980,3976,3972,3969,3965,3961,3958,3954,3950,3946,3942,3938,3934,3929,3925,3921,3917,3912,3908,3903,3899,3894,3889,3885,3880,3875,3870,3865,3861,3856,3851,3845,3840,3835,3830,3825,3819,3814,3808,3803,3797,3792,3786,3781,3775,3769,3763,3757,3751,3746,3740,3733,3727,3721,3715,3709,3703,3696,3690,3683,3677,3670,3664,3657,3651,3644,3637,3631,3624,3617,3610,3603,3596,3589,3582,3575,3568,3561,3553,3546,3539,3531,3524,3517,3509,3502,3494,3486,3479,3471,3463,3456,3448,3440,3432,3424,3416,3408,3400,3392,3384,3376,3368,3360,3351,3343,3335,3326,3318,3310,3301,3293,3284,3276,3267,3258,3250,3241,3232,3224,3215,3206,3197,3188,3179,3170,3161,3152,3143,3134,3125,3116,3107,3098,3089,3079,3070,3061,3051,3042,3033,3023,3014,3004,2995,2985,2976,2966,2957,2947,2937,2928,2918,2908,2899,2889,2879,2869,2859,2850,2840,2830,2820,2810,2800,2790,2780,2770,2760,2750,2740,2730,2720,2710,2699,2689,2679,2669,2659,2648,2638,2628,2618,2607,2597,2587,2576,2566,2556,2545,2535,2524,2514,2503,2493,2483,2472,2462,2451,2441,2430,2420,2409,2398,2388,2377,2367,2356,2346,2335,2324,2314,2303,2292,2282,2271,2260,2250,2239,2228,2218,2207,2196,2186,2175,2164,2154,2143,2132,2122,2111,2100,2089,2079,2068,2057,2047,2036,2025,2014,2004,1993,1982,1971,1961,1950,1939,1929,1918,1907,1897,1886,1875,1865,1854,1843,1833,1822,1811,1801,1790,1779,1769,1758,1747,1737,1726,1716,1705,1695,1684,1673,1663,1652,1642,1631,1621,1610,1600,1590,1579,1569,1558,1548,1537,1527,1517,1506,1496,1486,1475,1465,1455,1445,1434,1424,1414,1404,1394,1383,1373,1363,1353,1343,1333,1323,1313,1303,1293,1283,1273,1263,1253,1243,1234,1224,1214,1204,1194,1185,1175,1165,1156,1146,1136,1127,1117,1108,1098,1089,1079,1070,1060,1051,1042,1032,1023,1014,1004,995,986,977,968,959,950,941,932,923,914,905,896,887,878,869,861,852,843,835,826,817,809,800,792,783,775,767,758,750,742,733,725,717,709,701,693,685,677,669,661,653,645,637,630,622,614,607,599,591,584,576,569,562,554,547,540,532,525,518,511,504,497,490,483,476,469,462,456,449,442,436,429,423,416,410,403,397,390,384,378,372,366,360,353,347,342,336,330,324,318,312,307,301,296,290,285,279,274,268,263,258,253,248,242,237,232,228,223,218,213,208,204,199,194,190,185,181,176,172,168,164,159,155,151,147,143,139,135,132,128,124,121,117,113,110,106,103,100,96,93,90,87,84,81,78,75,72,69,67,64,61,59,56,54,51,49,46,44,42,40,38,36,34,32,30,28,26,25,23,21,20,18,17,16,14,13,12,11,10,9,8,7,6,5,4,4,3,2,2,1,1,1,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,3,4,4,5,6,7,8,9,10,11,12,13,14,16,17,18,20,21,23,25,26,28,30,32,34,36,38,40,42,44,46,49,51,54,56,59,61,64,67,69,72,75,78,81,84,87,90,93,96,100,103,106,110,113,117,121,124,128,132,135,139,143,147,151,155,159,164,168,172,176,181,185,190,194,199,204,208,213,218,223,228,232,237,242,248,253,258,263,268,274,279,285,290,296,301,307,312,318,324,330,336,342,347,353,360,366,372,378,384,390,397,403,410,416,423,429,436,442,449,456,462,469,476,483,490,497,504,511,518,525,532,540,547,554,562,569,576,584,591,599,607,614,622,630,637,645,653,661,669,677,685,693,701,709,717,725,733,742,750,758,767,775,783,792,800,809,817,826,835,843,852,861,869,878,887,896,905,914,923,932,941,950,959,968,977,986,995,1004,1014,1023,1032,1042,1051,1060,1070,1079,1089,1098,1108,1117,1127,1136,1146,1156,1165,1175,1185,1194,1204,1214,1224,1234,1243,1253,1263,1273,1283,1293,1303,1313,1323,1333,1343,1353,1363,1373,1383,1394,1404,1414,1424,1434,1445,1455,1465,1475,1486,1496,1506,1517,1527,1537,1548,1558,1569,1579,1590,1600,1610,1621,1631,1642,1652,1663,1673,1684,1695,1705,1716,1726,1737,1747,1758,1769,1779,1790,1801,1811,1822,1833,1843,1854,1865,1875,1886,1897,1907,1918,1929,1939,1950,1961,1971,1982,1993,2004,2014,2025,2036}; //loaded by python

    always @ (phase) begin
        //the phase is divided into two sections, where one set is an inversion of the other
        if (phase > SINE_RESOLUTION-1) begin
            signal <= -1 * sine_table[phase-SINE_RESOLUTION];
        end else begin
            signal <= sine_table[phase];
        end
    end
endmodule