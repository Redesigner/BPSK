`ifndef cross_comparison_sample_h
`define cross_comparison_sample_h
parameter signed [DATA_WIDTH-1:0] COMPARISON_TABLE [0:10*PREAMBLE_LENGTH - 1] = {0,1203,1946,1946,1203,0,-1203,-1946,-1946,-1203,0,1203,1946,1946,1203,0,-1203,-1946,-1946,-1203,0,1203,1946,1946,1203,0,-1203,-1946,-1946,-1203,0,1203,1946,1946,1203,0,-1203,-1946,-1946,-1203};
`endif