`ifndef preamble_params_h
`define preamble_params_h

localparam PREAMBLE_LENGTH = 4;
localparam PREAMBLE = 4'b1010;
localparam PREAMBLE_THRESHOLD = 79;

`endif