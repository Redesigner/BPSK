`ifndef cross_comparison_sample_h
`define cross_comparison_sample_h
parameter signed [DATA_WIDTH-1:0] COMPARISON_TABLE [0:$WAVELENGTH*PREAMBLE_LENGTH - 1] = $comparison_table;
`endif