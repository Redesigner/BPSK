`ifndef preamble_params_h
`define preamble_params_h

localparam PREAMBLE_LENGTH = $preamble_length;
localparam PREAMBLE = $preamble;
localparam PREAMBLE_THRESHOLD = $threshold;

`endif