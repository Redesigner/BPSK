`ifndef network_params_h
`define network_params_h

localparam NETWORK_WIDTH = 8;
localparam INDEX_WIDTH = 3;
localparam NETWORK_SLICES = 8;
localparam SORTING_WIDTH = NETWORK_SLICES * INDEX_WIDTH; 

`endif